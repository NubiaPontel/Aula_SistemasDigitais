/Trabalho, desenhar triângulos com verilog usando VGA/


module calc(
    input [10:0] p01x,
    input [10:0] p01y,
    input [10:0] p02x,
    input [10:0] p02y,
    input [10:0] p03x,
    input [10:0] p03y,
    output result
);

//result = (((p01.x - p03.x)*(p02.y - p03.y)) - ((p02.x - p03.x)*(p01.y - p03.y)));

wire signed [11:0] ss1;
wire signed [11:0] ss2;
wire signed [11:0] ss3;
wire signed [11:0] ss4;
wire signed [23:0] mm1;
wire signed [23:0] mm2;

assign s1 = p1x - p03x;
assign s2 = p2y - p03y;
assign s3 = p2x - p03x;
assign s4 = p1y - p03y;
assign m1 = s1 * ss2;
assign m2 = s3 * ss4;
assign result = mm1 > mm2;

endmodule

module videoMemoy(
	input wr,
	input [10:0] posx,
	input [10:0] posy,
	input [3:0] Redin,
	input [3:0] Greenin,
	input [3:0] Bluein,
	output [3:0] Redout,
	output [3:0] Greenout,
	output [3:0] Blueout
	);

	reg [11:0] mem [640:1][480:1];
	//307200 registradores de 12 bits ordenados em 640 linhas e 480 colunas.

	always @(posedge wr) begin
		if (wr == 1) begin
			mem[posx][posy][3:0] <= Red_in;
			mem[posx][posy][7:4] <= Green_in;
			mem[posx][posy][11:8] <= Blue_in;
		end
	end

	assign Red_out = mem[posx][posy][3:0];
	assign Green_out = mem[posx][posy][7:4];
	assign Blue_out = mem[posx][posy][11:8];

endmodule

module teste1;

reg clk = 0;
reg fim = 0;
reg wr;
reg [4:0] state = 0;
reg [10:0] posx;
reg [10:0] posy;
reg [4:0] triangulo;

reg [10:0] p01x;
reg [10:0] p01y;
reg [10:0] p02x;
reg [10:0] p02y;
reg [10:0] p03x;
reg [10:0] p03y;
reg [10:0] P0x;
reg [10:0] P0y;


reg [3:0] Red_in;
reg [3:0] Green_in;
reg [3:0] Blue_in;

wire [3:0] Red_out;
wire [3:0] Green_out;
wire [3:0] Blue_out;

wire t1, s1, s2, s3;

videoMemoy M(wr, pos_x, pos_y, Red_in, Green_in, Blue_in, Red_out, Green_out, Blue_out);

calc S1(p01x, p01y, p02x, p02y, p03x, p03y, t01);
calc S2(p01x, p01y, p02x, p02y, P0x, P0y, s01);
calc S3(p02x, p02y, p03x, p03y, P0x, P0y, s02);
calc S4(p03x, p03y, p01x, p01y, P0x, P0y, s03);

always #1 clk = ~clk;
always @(posedge clk) begin
	case(state)
	0: begin
		wr <= 0;
		pos_x <= 0;
		pos_y <= 0;
		triangulo <= 0;
		state <= 1;
	end
	1: begin
		p01x <= {$random} %639;
		p02x <= {$random} %639;
		p03x <= {$random} %639;
		p01y <= {$random} %479;
		p02y <= {$random} %479;
		p03y <= {$random} %479;

		P0x <= 0;
		P0y <= 0;
		triangulo <= triangulo + 1;
		state <= 2;
	end
	2: begin
		if (triangulo == 5) state <= 11;
		else begin
			if(P0x < 640) begin
				P0x <= P0x + 1;
				state <= 3;
			end
			else state <= 6;
		end
	end
	3: begin
		if(P0y < 480) begin
			P0y <= P0y + 1;
			state <= 4;
		end
		else begin
			Py <= 0;
			state <= 2;
		end
	end
	4: begin
		pos_x <= Px;
		pos_y <= Py;
		if (((t1 == s1) && (s1 == s2) && (s2 == s3))) begin
			case(triangulo)
			1: begin
				Red_in <= 4'b1111;
				Green_in <= 4'b0000;
				Blue_in <= 4'b0000;
			end
			2: begin
				Red_in <= 4'b0000;
				Green_in <= 4'b1111;
				Blue_in <= 4'b0000;
			end
			3: begin
				Red_in <= 4'b0000;
				Green_in <= 4'b0000;
				Blue_in <= 4'b1111;
			end
			4: begin
				Red_in <= 4'b1111;
				Green_in <= 4'b1111;
				Blue_in <= 4'b1111;
			end
			endcase
		end
		else begin
			Red_in <= 4'b0000;
			Green_in <= 4'b0000;
			Blue_in <= 4'b0000;
		end
		wr <= 1;
		state <= 5;
	end
	5: begin
		wr <= 0;
		state <= 3;
	end
	6: begin
		Px <= 0;
		Py <= 0;
		state <= 7;
	end
	7: begin
		if(Px < 640) begin
			Px <= Px + 1;
			state <= 8;
		end
		else state <= 1;
	end
	8: begin
		if(Py < 480) begin
			Py <= Py + 1;
			state <= 9;
		end
		else begin
			Py <= 0;
			state <= 7;
		end
	end
	9: begin
		pos_x <= Px;
		pos_y <= Py;
		state <= 10;
	end
	10: begin
		$display("\nTriangulo%d Mem[%d][%d] = R%d G%d B%d\n", triangulo, pos_x, pos_y, Red_out, Green_out, Blue_out);
		state <= 8;
	end
	11: $finish;
	endcase
end


endmodule
